// ********************************************************************
// >>>>>>>>>>>>>>>>>>>>>>>>> COPYRIGHT NOTICE <<<<<<<<<<<<<<<<<<<<<<<<<
// ********************************************************************
// File name    : segment.v
// Module name  : segment
// Author       : STEP
// Description  : segment initial
// Web          : www.stepfpga.com
// 
// --------------------------------------------------------------------
// Code Revision History : 
// --------------------------------------------------------------------
// Version: |Mod. Date:   |Changes Made:
// V1.0     |2017/03/02   |Initial ver
// --------------------------------------------------------------------
// Module Function:����ܵ�����ģ���ʼ��
 
module segment_LED (seg_data_1,seg_data_2,seg_led_1,seg_led_2);
 
	input [3:0] seg_data_1;						//�������Ҫ��ʾ0~9ʮ�����֣�����������Ҫ4λ����������
	input [3:0] seg_data_2;						//С��Ѿ�ϵڶ��������
	output [8:0] seg_led_1;						//��С��Ѿ�Ͽ���һ���������Ҫ9���ź� MSB~LSB=DIG��DP��G��F��E��D��C��B��A
	output [8:0] seg_led_2;						//��С��Ѿ�ϵڶ�������ܵĿ����ź�  MSB~LSB=DIG��DP��G��F��E��D��C��B��A
 
        reg [8:0] seg [15:0];                   //������һ��reg�͵�����������൱��һ��10*9�Ĵ洢�����洢��һ����10������ÿ������9λ��
 
        initial                                 //�ڹ��̿���ֻ�ܸ�reg�ͱ�����ֵ��Verilog�������ֹ��̿�always��initial
                                                //initial��always��ͬ���������ִֻ��һ��
	    begin
          seg[0] = 9'h3f;                       //�Դ洢���е�һ������ֵ9'b00_0011_1111,�൱�ڹ������ӵأ�DP���Ͳ�����7����ʾ����  0
	      seg[1] = 9'h06;                       //7����ʾ����  1
	      seg[2] = 9'h5b;                       //7����ʾ����  2
	      seg[3] = 9'h4f;                       //7����ʾ����  3
	      seg[4] = 9'h66;                       //7����ʾ����  4
	      seg[5] = 9'h6d;                       //7����ʾ����  5
	      seg[6] = 9'h7d;                       //7����ʾ����  6
	      seg[7] = 9'h07;                       //7����ʾ����  7
	      seg[8] = 9'h7f;                       //7����ʾ����  8
	      seg[9] = 9'h6f;                       //7����ʾ����  9
		  seg[10]= 9'hf7;						//	a
		  seg[11]= 9'h7c;	   					//  b
		  seg[12]= 9'h39;    					//  C           
		  seg[13]= 9'h5e;    					//  d
		  seg[14]= 9'h79;    					//  E
		  seg[15]= 9'h71;    					//  F
            end
 
        assign seg_led_1 = seg[seg_data_1];                         //������ֵ���������벻ͬ��λ��������������������9λ���
        assign seg_led_2 = seg[seg_data_2];
 
endmodule
